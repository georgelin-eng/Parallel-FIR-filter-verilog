// The FIR coefficients are generated at a sampling rate of 15000 kHz with a stop band of frequencies above 600 kHz

parameter width = 24;
parameter order = 53;

parameter integer FIRfilterCoeffs [order] = '{
    -3 ,
    -4 ,
    -5 ,
    -6 ,
    -8 ,
    -10 ,
    -11 ,
    -12 ,
    -12 ,
    -10 ,
    -6 ,
    0 ,
    9 ,
    22 ,
    38 ,
    57 ,
    79 ,
    104 ,
    130 ,
    157 ,
    183 ,
    208 ,
    230 ,
    248 ,
    262 ,
    270 ,
    273 ,
    270 ,
    262 ,
    248 ,
    230 ,
    208 ,
    183 ,
    157 ,
    130 ,
    104 ,
    79 ,
    57 ,
    38 ,
    22 ,
    9 ,
    0 ,
    -6 ,
    -10 ,
    -12 ,
    -12 ,
    -11 ,
    -10 ,
    -8 ,
    -6 ,
    -5 ,
    -4 ,
    -3};