
/* ----------------------------
* 
* Author:  George Lin
* Purpose: Composed of generator, driver, interface, monitor, and scoreboard to 
*          increase modularity and scalability of testing environment. 
* 
* 
-----------------------------  */

module FIR_testBench_TOP();
// instantiation of the DUT


endmodule


class FIR_item
    // transaction object

    
endclass

class FIR_interface
endclass

class generator
endclass

class driver
endclass


class monitor
    
endclass

class scoreboard


endclass

class env
    driver      d0;
    monitor     m0;
    generator   g0;
    scoreboard  s0;


    

endclass

class test
endclass
